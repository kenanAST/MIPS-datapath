module and2(d, b, c); 
    input d, b;
    output c;     
    assign c = d & b; 
endmodule 